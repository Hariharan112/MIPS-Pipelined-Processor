//mips control module only for ORI,LW,SUB, XOr